
parameter I2C_ADDR_WIDTH = 7;
parameter I2C_DATA_WIDTH = 8;

//typedef enum bit {WRITE = 0, READ =1} i2c_op_t;