package defines_pkg;

typedef enum bit {WRITE = 0, READ =1} i2c_op_t;

endpackage